library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

library work;

entity test2 is
	port(
		test_i	: in std_logic
	);
end test2;

architecture rtl of test2 is
begin
end rtl;
