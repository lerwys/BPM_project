library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

library work;

entity test is
	port(
		test_i	: in std_logic
	);
end test;

architecture rtl of test is
begin
end rtl;
